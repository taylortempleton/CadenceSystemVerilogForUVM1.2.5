/*-----------------------------------------------------------------
From the Cadence "Essential SystemVerilog for UVM" training course
Copyright Cadence Design Systems (c)2019

2022 Jan 18
taylor.templeton@gmail.com
Solution to lab04
-----------------------------------------------------------------*/

package packet_pkg;
 
`include "packet_data.sv" 

endpackage