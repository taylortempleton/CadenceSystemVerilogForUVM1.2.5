/*-----------------------------------------------------------------
From the Cadence "Essential SystemVerilog for UVM" training course
Copyright Cadence Design Systems (c)2019

2022 Jan 18
taylor.templeton@gmail.com
Solution to lab05
-----------------------------------------------------------------*/

package packet_pkg;
 
`include "packet_data.sv" 
`include "component_base.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "packet_vc.sv"

endpackage